library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

--hazard entity for dependency in arithmetic and logical instructions
entity hazard_EX is
	port( RREX_opcode, EXMA_opcode, MAWB_opcode: in std_logic_vector(3 downto 0); 
		  RREX_11_9, RREX_8_6, EXMA_11_9, MAWB_11_9, MAWB_8_6, MAWB_5_3: in std_logic_vector(2 downto 0);
          EXMA_1_0, MAWB_1_0, EXMA_flags, MAWB_flags : in std_logic_vector(1 downto 0);
		  disable_IFID, disable_IDRR, disable_RREX: out std_logic;
          alu2a_mux, alu2b_mux, PC_mux : out std_logic_vector(2 downto 0));  -- disable means we don't write anything in pipelined register in WB stage
end entity;

architecture hazardous of hazard_EX is
signal jalr_jri_jal , beq,ble,blt, add_nand__load_op :  std_logic := '0';
begin
add_nand__load_op <= '1' when(
    ((EXMA_opcode = "0001" or EXMA_opcode = "0010") and EXMA_1_0 = "00") or
    ((EXMA_opcode = "0001" or EXMA_opcode = "0010") and EXMA_1_0 = "10" and EXMA_flags(1 downto 1) = '1') or
    ((EXMA_opcode = "0001" or EXMA_opcode = "0010") and EXMA_1_0 = "01" and EXMA_flags(0 downto 0) = '1') or
    ((EXMA_opcode = "0001" or EXMA_opcode = "0010") and EXMA_1_0 = "11" and EXMA_flags(1 downto 0) = "11") or
    ((MAWB_opcode = "0001" or MAWB_opcode = "0010") and MAWB_1_0 = "00") or
    ((MAWB_opcode = "0001" or MAWB_opcode = "0010") and MAWB_1_0 = "10" and MAWB_flags(1 downto 1) = '1') or
    ((MAWB_opcode = "0001" or MAWB_opcode = "0010") and MAWB_1_0 = "01" and MAWB_flags(0 downto 0) = '1') or
    ((MAWB_opcode = "0001" or MAWB_opcode = "0010") and MAWB_1_0 = "11" and MAWB_flags(1 downto 0) = "11") or
    (EXMA_opcode = "0000") or (MAWB_opcode = "0000") or 
    (EXMA_opcode = "0011" or EXMA_opcode = "0100") or
    (MAWB_opcode = "0011" or MAWB_opcode = "0100")
) else '0';
--PC_mux (8x1 16 bit) if S= 010 => ALU4 , 001 =>ALU2 , 000 =>ALU1 011 => SE7 100 => Mem2D
PC_mux <=   "001" when(((EXMA_5_3 = "000" and (EXMA_opcode = "0001" or EXMA_opcode = "0010") ) or --all conditional A/L
                        (EXMA_opcode = "0000" and EXMA_8_6 ="000" )) and add_nand__load_op) else
            "010" when((EXMA_opcode = "1100" or "1101" or "1111") or (EXMA_opcode = "1000"  and (EXMA_flags = '01')) or      --all branch +jump
                       (EXMA_opcode = "1000"  and (EXMA_flags = '10')) or (EXMA_opcode = "1001"  and (EXMA_flags = '10' or '11'))) else
            "011" when (EXMA_11_9 = "000" and EXMA_opcode = "0011" and add_nand__load_op) else   --LLI
            "100" when (MAWB_11_9 = "000" and  MAWB_opcode = "0100" and add_nand__load_op)   --LW 
    else    "000";

-- alu2
alu2a_haz_mux <= "001" when(((RREX_11_9 = EXMA_5_3 and (EXMA_opcode = "0001" or EXMA_opcode = "0010")) or ((RREX_11_9 = EXMA_8_6) and EXMA_opcode = "0000")) and alu_nand_op) else
                 "010" when(((RREX_11_9 = MAWB_5_3 and (MAWB_opcode = "0001" or MAWB_opcode = "0010")) or ((RREX_11_9 = MAWB_8_6) and MAWB_opcode = "0000"))  and alu_nand_op) else
                 "011" when(RREX_11_9 = EXMA_11_9 and EXMA_opcode = "0011" and add_nand__load_op) else
                 "100" when(RREX_11_9 = MAWB_11_9 and MAWB_opcode = "0100" and add_nand__load_op) else
                 "000"
alu2b_haz_mux <= "001" when(((RREX_8_6 = EXMA_5_3 and (EXMA_opcode = "0001" or EXMA_opcode = "0010")) or ((RREX_8_6 = EXMA_8_6) and EXMA_opcode = "0000")) and alu_nand_op) else;
                 "010" when(((RREX_8_6 = MAWB_5_3 and (MAWB_opcode = "0001" or MAWB_opcode = "0010")) or ((RREX_8_6 = MAWB_8_6) and MAWB_opcode = "0000")) and alu_nand_op) else
                 "011" when(RREX_8_6 = EXMA_11_9 and EXMA_opcode = "0011" and add_nand__load_op) else
                 "100" when(RREX_8_6 = MAWB_11_9 and MAWB_opcode = "0100" and add_nand__load_op) else
                 "000"


jalr_jri_jal <= '1' when(RREX_opcode = "1100" or "1101" or "1111") else '0'; -- basically when there is all unconditional jump statements jal,jlr,jri then disable if_id,id_rr,rr_ex in nxt clk cycle
beq <= '1' when(RREX_opcode = "1000"  and (EXMA_flags = "01")) else '0';
blt <= '1' when(RREX_opcode = "1000"  and (EXMA_flags = "10")) else '0';
ble <= '1' when(RREX_opcode = "1001"  and (EXMA_flags = "10" or '11')) else '0';  -- correct vedika's alu

 disable_IFID <= '1'  when(jalr_jri_jal='1' or beq='1' or ble='1' or blt='1' or (PC_mux = "01" or PC_mux = "10"));
 disable_IDRR <= '1' when (jalr_jri_jal='1' or beq='1' or ble='1' or blt='1' or (PC_mux = "01" or PC_mux = "10"));
 disable_RREX <= '1' when (jalr_jri_jal or beq or ble or blt or (PC_mux = "01" or PC_mux = "10"));

 -- need to make rf_w, mem2_w, flag_w =0
end architecture;
